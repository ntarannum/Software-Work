// slave.v

// Generated using ACDS version 13.1 162 at 2018.11.27.10:02:01

`timescale 1 ps / 1 ps
module slave (
		input  wire       clk_clk,              //           clk.clk
		output wire [1:0] et_led1_export,       //       et_led1.export
		output wire [1:0] et_led2_export,       //       et_led2.export
		input  wire       spi_0_MISO,           //         spi_0.MISO
		output wire       spi_0_MOSI,           //              .MOSI
		output wire       spi_0_SCLK,           //              .SCLK
		output wire       spi_0_SS_n,           //              .SS_n
		input  wire       spi_can_int_n_export, // spi_can_int_n.export
		input  wire       et_pb_1_export,       //       et_pb_1.export
		input  wire       et_pb_2_export,       //       et_pb_2.export
		output wire [3:0] tt_led_export,        //        tt_led.export
		input  wire       tt_pb_1_export,       //       tt_pb_1.export
		output wire       tt_test_export        //       tt_test.export
	);

	wire  [31:0] mm_interconnect_0_et_leds2_s1_writedata;                     // mm_interconnect_0:et_leds2_s1_writedata -> et_leds2:writedata
	wire   [1:0] mm_interconnect_0_et_leds2_s1_address;                       // mm_interconnect_0:et_leds2_s1_address -> et_leds2:address
	wire         mm_interconnect_0_et_leds2_s1_chipselect;                    // mm_interconnect_0:et_leds2_s1_chipselect -> et_leds2:chipselect
	wire         mm_interconnect_0_et_leds2_s1_write;                         // mm_interconnect_0:et_leds2_s1_write -> et_leds2:write_n
	wire  [31:0] mm_interconnect_0_et_leds2_s1_readdata;                      // et_leds2:readdata -> mm_interconnect_0:et_leds2_s1_readdata
	wire  [31:0] mm_interconnect_0_msg_buf_mutex_s1_writedata;                // mm_interconnect_0:msg_buf_mutex_s1_writedata -> msg_buf_mutex:data_from_cpu
	wire   [0:0] mm_interconnect_0_msg_buf_mutex_s1_address;                  // mm_interconnect_0:msg_buf_mutex_s1_address -> msg_buf_mutex:address
	wire         mm_interconnect_0_msg_buf_mutex_s1_chipselect;               // mm_interconnect_0:msg_buf_mutex_s1_chipselect -> msg_buf_mutex:chipselect
	wire         mm_interconnect_0_msg_buf_mutex_s1_write;                    // mm_interconnect_0:msg_buf_mutex_s1_write -> msg_buf_mutex:write
	wire         mm_interconnect_0_msg_buf_mutex_s1_read;                     // mm_interconnect_0:msg_buf_mutex_s1_read -> msg_buf_mutex:read
	wire  [31:0] mm_interconnect_0_msg_buf_mutex_s1_readdata;                 // msg_buf_mutex:data_to_cpu -> mm_interconnect_0:msg_buf_mutex_s1_readdata
	wire  [15:0] mm_interconnect_0_et_spi_0_spi_control_port_writedata;       // mm_interconnect_0:et_spi_0_spi_control_port_writedata -> et_spi_0:data_from_cpu
	wire   [2:0] mm_interconnect_0_et_spi_0_spi_control_port_address;         // mm_interconnect_0:et_spi_0_spi_control_port_address -> et_spi_0:mem_addr
	wire         mm_interconnect_0_et_spi_0_spi_control_port_chipselect;      // mm_interconnect_0:et_spi_0_spi_control_port_chipselect -> et_spi_0:spi_select
	wire         mm_interconnect_0_et_spi_0_spi_control_port_write;           // mm_interconnect_0:et_spi_0_spi_control_port_write -> et_spi_0:write_n
	wire         mm_interconnect_0_et_spi_0_spi_control_port_read;            // mm_interconnect_0:et_spi_0_spi_control_port_read -> et_spi_0:read_n
	wire  [15:0] mm_interconnect_0_et_spi_0_spi_control_port_readdata;        // et_spi_0:data_to_cpu -> mm_interconnect_0:et_spi_0_spi_control_port_readdata
	wire  [31:0] mm_interconnect_0_et_core_memory_s1_writedata;               // mm_interconnect_0:ET_Core_Memory_s1_writedata -> ET_Core_Memory:writedata
	wire  [11:0] mm_interconnect_0_et_core_memory_s1_address;                 // mm_interconnect_0:ET_Core_Memory_s1_address -> ET_Core_Memory:address
	wire         mm_interconnect_0_et_core_memory_s1_chipselect;              // mm_interconnect_0:ET_Core_Memory_s1_chipselect -> ET_Core_Memory:chipselect
	wire         mm_interconnect_0_et_core_memory_s1_clken;                   // mm_interconnect_0:ET_Core_Memory_s1_clken -> ET_Core_Memory:clken
	wire         mm_interconnect_0_et_core_memory_s1_write;                   // mm_interconnect_0:ET_Core_Memory_s1_write -> ET_Core_Memory:write
	wire  [31:0] mm_interconnect_0_et_core_memory_s1_readdata;                // ET_Core_Memory:readdata -> mm_interconnect_0:ET_Core_Memory_s1_readdata
	wire   [3:0] mm_interconnect_0_et_core_memory_s1_byteenable;              // mm_interconnect_0:ET_Core_Memory_s1_byteenable -> ET_Core_Memory:byteenable
	wire  [15:0] mm_interconnect_0_tt_timer_1_s1_writedata;                   // mm_interconnect_0:tt_timer_1_s1_writedata -> tt_timer_1:writedata
	wire   [2:0] mm_interconnect_0_tt_timer_1_s1_address;                     // mm_interconnect_0:tt_timer_1_s1_address -> tt_timer_1:address
	wire         mm_interconnect_0_tt_timer_1_s1_chipselect;                  // mm_interconnect_0:tt_timer_1_s1_chipselect -> tt_timer_1:chipselect
	wire         mm_interconnect_0_tt_timer_1_s1_write;                       // mm_interconnect_0:tt_timer_1_s1_write -> tt_timer_1:write_n
	wire  [15:0] mm_interconnect_0_tt_timer_1_s1_readdata;                    // tt_timer_1:readdata -> mm_interconnect_0:tt_timer_1_s1_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire  [31:0] mm_interconnect_0_tt_core_memory_s1_writedata;               // mm_interconnect_0:TT_core_memory_s1_writedata -> TT_core_memory:writedata
	wire  [11:0] mm_interconnect_0_tt_core_memory_s1_address;                 // mm_interconnect_0:TT_core_memory_s1_address -> TT_core_memory:address
	wire         mm_interconnect_0_tt_core_memory_s1_chipselect;              // mm_interconnect_0:TT_core_memory_s1_chipselect -> TT_core_memory:chipselect
	wire         mm_interconnect_0_tt_core_memory_s1_clken;                   // mm_interconnect_0:TT_core_memory_s1_clken -> TT_core_memory:clken
	wire         mm_interconnect_0_tt_core_memory_s1_write;                   // mm_interconnect_0:TT_core_memory_s1_write -> TT_core_memory:write
	wire  [31:0] mm_interconnect_0_tt_core_memory_s1_readdata;                // TT_core_memory:readdata -> mm_interconnect_0:TT_core_memory_s1_readdata
	wire   [3:0] mm_interconnect_0_tt_core_memory_s1_byteenable;              // mm_interconnect_0:TT_core_memory_s1_byteenable -> TT_core_memory:byteenable
	wire   [1:0] mm_interconnect_0_et_pb_2_s1_address;                        // mm_interconnect_0:et_pb_2_s1_address -> et_pb_2:address
	wire  [31:0] mm_interconnect_0_et_pb_2_s1_readdata;                       // et_pb_2:readdata -> mm_interconnect_0:et_pb_2_s1_readdata
	wire  [31:0] mm_interconnect_0_et_leds1_s1_writedata;                     // mm_interconnect_0:et_leds1_s1_writedata -> et_leds1:writedata
	wire   [1:0] mm_interconnect_0_et_leds1_s1_address;                       // mm_interconnect_0:et_leds1_s1_address -> et_leds1:address
	wire         mm_interconnect_0_et_leds1_s1_chipselect;                    // mm_interconnect_0:et_leds1_s1_chipselect -> et_leds1:chipselect
	wire         mm_interconnect_0_et_leds1_s1_write;                         // mm_interconnect_0:et_leds1_s1_write -> et_leds1:write_n
	wire  [31:0] mm_interconnect_0_et_leds1_s1_readdata;                      // et_leds1:readdata -> mm_interconnect_0:et_leds1_s1_readdata
	wire  [31:0] mm_interconnect_0_msg_buf_ram_s1_writedata;                  // mm_interconnect_0:msg_buf_ram_s1_writedata -> msg_buf_ram:writedata
	wire   [7:0] mm_interconnect_0_msg_buf_ram_s1_address;                    // mm_interconnect_0:msg_buf_ram_s1_address -> msg_buf_ram:address
	wire         mm_interconnect_0_msg_buf_ram_s1_chipselect;                 // mm_interconnect_0:msg_buf_ram_s1_chipselect -> msg_buf_ram:chipselect
	wire         mm_interconnect_0_msg_buf_ram_s1_clken;                      // mm_interconnect_0:msg_buf_ram_s1_clken -> msg_buf_ram:clken
	wire         mm_interconnect_0_msg_buf_ram_s1_write;                      // mm_interconnect_0:msg_buf_ram_s1_write -> msg_buf_ram:write
	wire  [31:0] mm_interconnect_0_msg_buf_ram_s1_readdata;                   // msg_buf_ram:readdata -> mm_interconnect_0:msg_buf_ram_s1_readdata
	wire   [3:0] mm_interconnect_0_msg_buf_ram_s1_byteenable;                 // mm_interconnect_0:msg_buf_ram_s1_byteenable -> msg_buf_ram:byteenable
	wire   [1:0] mm_interconnect_0_tt_pb_1_s1_address;                        // mm_interconnect_0:tt_pb_1_s1_address -> tt_pb_1:address
	wire  [31:0] mm_interconnect_0_tt_pb_1_s1_readdata;                       // tt_pb_1:readdata -> mm_interconnect_0:tt_pb_1_s1_readdata
	wire         et_core_data_master_waitrequest;                             // mm_interconnect_0:ET_Core_data_master_waitrequest -> ET_Core:d_waitrequest
	wire  [31:0] et_core_data_master_writedata;                               // ET_Core:d_writedata -> mm_interconnect_0:ET_Core_data_master_writedata
	wire  [15:0] et_core_data_master_address;                                 // ET_Core:d_address -> mm_interconnect_0:ET_Core_data_master_address
	wire         et_core_data_master_write;                                   // ET_Core:d_write -> mm_interconnect_0:ET_Core_data_master_write
	wire         et_core_data_master_read;                                    // ET_Core:d_read -> mm_interconnect_0:ET_Core_data_master_read
	wire  [31:0] et_core_data_master_readdata;                                // mm_interconnect_0:ET_Core_data_master_readdata -> ET_Core:d_readdata
	wire         et_core_data_master_debugaccess;                             // ET_Core:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:ET_Core_data_master_debugaccess
	wire   [3:0] et_core_data_master_byteenable;                              // ET_Core:d_byteenable -> mm_interconnect_0:ET_Core_data_master_byteenable
	wire         mm_interconnect_0_tt_core_jtag_debug_module_waitrequest;     // TT_Core:jtag_debug_module_waitrequest -> mm_interconnect_0:TT_Core_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_tt_core_jtag_debug_module_writedata;       // mm_interconnect_0:TT_Core_jtag_debug_module_writedata -> TT_Core:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_tt_core_jtag_debug_module_address;         // mm_interconnect_0:TT_Core_jtag_debug_module_address -> TT_Core:jtag_debug_module_address
	wire         mm_interconnect_0_tt_core_jtag_debug_module_write;           // mm_interconnect_0:TT_Core_jtag_debug_module_write -> TT_Core:jtag_debug_module_write
	wire         mm_interconnect_0_tt_core_jtag_debug_module_read;            // mm_interconnect_0:TT_Core_jtag_debug_module_read -> TT_Core:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_tt_core_jtag_debug_module_readdata;        // TT_Core:jtag_debug_module_readdata -> mm_interconnect_0:TT_Core_jtag_debug_module_readdata
	wire         mm_interconnect_0_tt_core_jtag_debug_module_debugaccess;     // mm_interconnect_0:TT_Core_jtag_debug_module_debugaccess -> TT_Core:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_tt_core_jtag_debug_module_byteenable;      // mm_interconnect_0:TT_Core_jtag_debug_module_byteenable -> TT_Core:jtag_debug_module_byteenable
	wire         et_core_instruction_master_waitrequest;                      // mm_interconnect_0:ET_Core_instruction_master_waitrequest -> ET_Core:i_waitrequest
	wire  [15:0] et_core_instruction_master_address;                          // ET_Core:i_address -> mm_interconnect_0:ET_Core_instruction_master_address
	wire         et_core_instruction_master_read;                             // ET_Core:i_read -> mm_interconnect_0:ET_Core_instruction_master_read
	wire  [31:0] et_core_instruction_master_readdata;                         // mm_interconnect_0:ET_Core_instruction_master_readdata -> ET_Core:i_readdata
	wire         mm_interconnect_0_et_core_jtag_debug_module_waitrequest;     // ET_Core:jtag_debug_module_waitrequest -> mm_interconnect_0:ET_Core_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_et_core_jtag_debug_module_writedata;       // mm_interconnect_0:ET_Core_jtag_debug_module_writedata -> ET_Core:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_et_core_jtag_debug_module_address;         // mm_interconnect_0:ET_Core_jtag_debug_module_address -> ET_Core:jtag_debug_module_address
	wire         mm_interconnect_0_et_core_jtag_debug_module_write;           // mm_interconnect_0:ET_Core_jtag_debug_module_write -> ET_Core:jtag_debug_module_write
	wire         mm_interconnect_0_et_core_jtag_debug_module_read;            // mm_interconnect_0:ET_Core_jtag_debug_module_read -> ET_Core:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_et_core_jtag_debug_module_readdata;        // ET_Core:jtag_debug_module_readdata -> mm_interconnect_0:ET_Core_jtag_debug_module_readdata
	wire         mm_interconnect_0_et_core_jtag_debug_module_debugaccess;     // mm_interconnect_0:ET_Core_jtag_debug_module_debugaccess -> ET_Core:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_et_core_jtag_debug_module_byteenable;      // mm_interconnect_0:ET_Core_jtag_debug_module_byteenable -> ET_Core:jtag_debug_module_byteenable
	wire  [31:0] mm_interconnect_0_et_spican_int_s1_writedata;                // mm_interconnect_0:et_spican_int_s1_writedata -> et_spican_int:writedata
	wire   [1:0] mm_interconnect_0_et_spican_int_s1_address;                  // mm_interconnect_0:et_spican_int_s1_address -> et_spican_int:address
	wire         mm_interconnect_0_et_spican_int_s1_chipselect;               // mm_interconnect_0:et_spican_int_s1_chipselect -> et_spican_int:chipselect
	wire         mm_interconnect_0_et_spican_int_s1_write;                    // mm_interconnect_0:et_spican_int_s1_write -> et_spican_int:write_n
	wire  [31:0] mm_interconnect_0_et_spican_int_s1_readdata;                 // et_spican_int:readdata -> mm_interconnect_0:et_spican_int_s1_readdata
	wire  [31:0] mm_interconnect_0_tt_leds_s1_writedata;                      // mm_interconnect_0:tt_leds_s1_writedata -> tt_leds:writedata
	wire   [1:0] mm_interconnect_0_tt_leds_s1_address;                        // mm_interconnect_0:tt_leds_s1_address -> tt_leds:address
	wire         mm_interconnect_0_tt_leds_s1_chipselect;                     // mm_interconnect_0:tt_leds_s1_chipselect -> tt_leds:chipselect
	wire         mm_interconnect_0_tt_leds_s1_write;                          // mm_interconnect_0:tt_leds_s1_write -> tt_leds:write_n
	wire  [31:0] mm_interconnect_0_tt_leds_s1_readdata;                       // tt_leds:readdata -> mm_interconnect_0:tt_leds_s1_readdata
	wire         tt_core_data_master_waitrequest;                             // mm_interconnect_0:TT_Core_data_master_waitrequest -> TT_Core:d_waitrequest
	wire  [31:0] tt_core_data_master_writedata;                               // TT_Core:d_writedata -> mm_interconnect_0:TT_Core_data_master_writedata
	wire  [15:0] tt_core_data_master_address;                                 // TT_Core:d_address -> mm_interconnect_0:TT_Core_data_master_address
	wire         tt_core_data_master_write;                                   // TT_Core:d_write -> mm_interconnect_0:TT_Core_data_master_write
	wire         tt_core_data_master_read;                                    // TT_Core:d_read -> mm_interconnect_0:TT_Core_data_master_read
	wire  [31:0] tt_core_data_master_readdata;                                // mm_interconnect_0:TT_Core_data_master_readdata -> TT_Core:d_readdata
	wire         tt_core_data_master_debugaccess;                             // TT_Core:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:TT_Core_data_master_debugaccess
	wire   [3:0] tt_core_data_master_byteenable;                              // TT_Core:d_byteenable -> mm_interconnect_0:TT_Core_data_master_byteenable
	wire   [1:0] mm_interconnect_0_et_pb_1_s1_address;                        // mm_interconnect_0:et_pb_1_s1_address -> et_pb_1:address
	wire  [31:0] mm_interconnect_0_et_pb_1_s1_readdata;                       // et_pb_1:readdata -> mm_interconnect_0:et_pb_1_s1_readdata
	wire  [31:0] mm_interconnect_0_pio_0_s1_writedata;                        // mm_interconnect_0:pio_0_s1_writedata -> pio_0:writedata
	wire   [1:0] mm_interconnect_0_pio_0_s1_address;                          // mm_interconnect_0:pio_0_s1_address -> pio_0:address
	wire         mm_interconnect_0_pio_0_s1_chipselect;                       // mm_interconnect_0:pio_0_s1_chipselect -> pio_0:chipselect
	wire         mm_interconnect_0_pio_0_s1_write;                            // mm_interconnect_0:pio_0_s1_write -> pio_0:write_n
	wire  [31:0] mm_interconnect_0_pio_0_s1_readdata;                         // pio_0:readdata -> mm_interconnect_0:pio_0_s1_readdata
	wire         tt_core_instruction_master_waitrequest;                      // mm_interconnect_0:TT_Core_instruction_master_waitrequest -> TT_Core:i_waitrequest
	wire  [15:0] tt_core_instruction_master_address;                          // TT_Core:i_address -> mm_interconnect_0:TT_Core_instruction_master_address
	wire         tt_core_instruction_master_read;                             // TT_Core:i_read -> mm_interconnect_0:TT_Core_instruction_master_read
	wire  [31:0] tt_core_instruction_master_readdata;                         // mm_interconnect_0:TT_Core_instruction_master_readdata -> TT_Core:i_readdata
	wire         irq_mapper_receiver0_irq;                                    // et_spi_0:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                    // et_spican_int:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver2_irq
	wire  [31:0] et_core_d_irq_irq;                                           // irq_mapper:sender_irq -> ET_Core:d_irq
	wire         irq_mapper_001_receiver0_irq;                                // tt_timer_1:irq -> irq_mapper_001:receiver0_irq
	wire  [31:0] tt_core_d_irq_irq;                                           // irq_mapper_001:sender_irq -> TT_Core:d_irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> rst_controller_001:reset_in0
	wire         tt_core_jtag_debug_module_reset_reset;                       // TT_Core:jtag_debug_module_resetrequest -> [rst_controller:reset_in0, rst_controller_001:reset_in2]
	wire         et_core_jtag_debug_module_reset_reset;                       // ET_Core:jtag_debug_module_resetrequest -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	wire         rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [ET_Core:reset_n, ET_Core_Memory:reset, TT_Core:reset_n, TT_core_memory:reset, et_leds1:reset_n, et_leds2:reset_n, et_pb_1:reset_n, et_pb_2:reset_n, et_spi_0:reset_n, et_spican_int:reset_n, irq_mapper:reset, irq_mapper_001:reset, jtag_uart_0:rst_n, mm_interconnect_0:ET_Core_reset_n_reset_bridge_in_reset_reset, msg_buf_mutex:reset_n, msg_buf_ram:reset, pio_0:reset_n, rst_translator:in_reset, tt_leds:reset_n, tt_pb_1:reset_n, tt_timer_1:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                      // rst_controller_001:reset_req -> [ET_Core:reset_req, ET_Core_Memory:reset_req, TT_Core:reset_req, TT_core_memory:reset_req, msg_buf_ram:reset_req, rst_translator:reset_req_in]

	slave_ET_Core et_core (
		.clk                                   (clk_clk),                                                 //                       clk.clk
		.reset_n                               (~rst_controller_001_reset_out_reset),                     //                   reset_n.reset_n
		.reset_req                             (rst_controller_001_reset_out_reset_req),                  //                          .reset_req
		.d_address                             (et_core_data_master_address),                             //               data_master.address
		.d_byteenable                          (et_core_data_master_byteenable),                          //                          .byteenable
		.d_read                                (et_core_data_master_read),                                //                          .read
		.d_readdata                            (et_core_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (et_core_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (et_core_data_master_write),                               //                          .write
		.d_writedata                           (et_core_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (et_core_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (et_core_instruction_master_address),                      //        instruction_master.address
		.i_read                                (et_core_instruction_master_read),                         //                          .read
		.i_readdata                            (et_core_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (et_core_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (et_core_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (et_core_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_et_core_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_et_core_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_et_core_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_et_core_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_et_core_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_et_core_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_et_core_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_et_core_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                         // custom_instruction_master.readra
	);

	slave_ET_Core_Memory et_core_memory (
		.clk        (clk_clk),                                        //   clk1.clk
		.address    (mm_interconnect_0_et_core_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_et_core_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_et_core_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_et_core_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_et_core_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_et_core_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_et_core_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req)          //       .reset_req
	);

	slave_et_leds1 et_leds1 (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_et_leds1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_et_leds1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_et_leds1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_et_leds1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_et_leds1_s1_readdata),   //                    .readdata
		.out_port   (et_led1_export)                            // external_connection.export
	);

	slave_et_leds1 et_leds2 (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_et_leds2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_et_leds2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_et_leds2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_et_leds2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_et_leds2_s1_readdata),   //                    .readdata
		.out_port   (et_led2_export)                            // external_connection.export
	);

	slave_et_spi_0 et_spi_0 (
		.clk           (clk_clk),                                                //              clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),                    //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_et_spi_0_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_et_spi_0_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_et_spi_0_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_et_spi_0_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_et_spi_0_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_et_spi_0_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver0_irq),                               //              irq.irq
		.MISO          (spi_0_MISO),                                             //         external.export
		.MOSI          (spi_0_MOSI),                                             //                 .export
		.SCLK          (spi_0_SCLK),                                             //                 .export
		.SS_n          (spi_0_SS_n)                                              //                 .export
	);

	slave_et_spican_int et_spican_int (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_et_spican_int_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_et_spican_int_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_et_spican_int_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_et_spican_int_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_et_spican_int_s1_readdata),   //                    .readdata
		.in_port    (spi_can_int_n_export),                          // external_connection.export
		.irq        (irq_mapper_receiver1_irq)                       //                 irq.irq
	);

	slave_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                         //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver2_irq)                                     //               irq.irq
	);

	slave_et_pb_1 et_pb_1 (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),   //               reset.reset_n
		.address  (mm_interconnect_0_et_pb_1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_et_pb_1_s1_readdata), //                    .readdata
		.in_port  (et_pb_1_export)                         // external_connection.export
	);

	slave_et_pb_1 et_pb_2 (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),   //               reset.reset_n
		.address  (mm_interconnect_0_et_pb_2_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_et_pb_2_s1_readdata), //                    .readdata
		.in_port  (et_pb_2_export)                         // external_connection.export
	);

	slave_TT_Core tt_core (
		.clk                                   (clk_clk),                                                 //                       clk.clk
		.reset_n                               (~rst_controller_001_reset_out_reset),                     //                   reset_n.reset_n
		.reset_req                             (rst_controller_001_reset_out_reset_req),                  //                          .reset_req
		.d_address                             (tt_core_data_master_address),                             //               data_master.address
		.d_byteenable                          (tt_core_data_master_byteenable),                          //                          .byteenable
		.d_read                                (tt_core_data_master_read),                                //                          .read
		.d_readdata                            (tt_core_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (tt_core_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (tt_core_data_master_write),                               //                          .write
		.d_writedata                           (tt_core_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (tt_core_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (tt_core_instruction_master_address),                      //        instruction_master.address
		.i_read                                (tt_core_instruction_master_read),                         //                          .read
		.i_readdata                            (tt_core_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (tt_core_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (tt_core_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (tt_core_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_tt_core_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_tt_core_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_tt_core_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_tt_core_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_tt_core_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_tt_core_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_tt_core_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_tt_core_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                         // custom_instruction_master.readra
	);

	slave_TT_core_memory tt_core_memory (
		.clk        (clk_clk),                                        //   clk1.clk
		.address    (mm_interconnect_0_tt_core_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_tt_core_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_tt_core_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_tt_core_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_tt_core_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_tt_core_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_tt_core_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req)          //       .reset_req
	);

	slave_tt_leds tt_leds (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_tt_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_tt_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_tt_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_tt_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_tt_leds_s1_readdata),   //                    .readdata
		.out_port   (tt_led_export)                            // external_connection.export
	);

	slave_et_pb_1 tt_pb_1 (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),   //               reset.reset_n
		.address  (mm_interconnect_0_tt_pb_1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_tt_pb_1_s1_readdata), //                    .readdata
		.in_port  (tt_pb_1_export)                         // external_connection.export
	);

	slave_msg_buf_mutex msg_buf_mutex (
		.reset_n       (~rst_controller_001_reset_out_reset),           // reset.reset_n
		.clk           (clk_clk),                                       //   clk.clk
		.chipselect    (mm_interconnect_0_msg_buf_mutex_s1_chipselect), //    s1.chipselect
		.data_from_cpu (mm_interconnect_0_msg_buf_mutex_s1_writedata),  //      .writedata
		.read          (mm_interconnect_0_msg_buf_mutex_s1_read),       //      .read
		.write         (mm_interconnect_0_msg_buf_mutex_s1_write),      //      .write
		.data_to_cpu   (mm_interconnect_0_msg_buf_mutex_s1_readdata),   //      .readdata
		.address       (mm_interconnect_0_msg_buf_mutex_s1_address)     //      .address
	);

	slave_msg_buf_ram msg_buf_ram (
		.clk        (clk_clk),                                     //   clk1.clk
		.address    (mm_interconnect_0_msg_buf_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_msg_buf_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_msg_buf_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_msg_buf_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_msg_buf_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_msg_buf_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_msg_buf_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),          // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req)       //       .reset_req
	);

	slave_pio_0 pio_0 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),   //               reset.reset_n
		.address    (mm_interconnect_0_pio_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_0_s1_readdata),   //                    .readdata
		.out_port   (tt_test_export)                         // external_connection.export
	);

	slave_tt_timer_1 tt_timer_1 (
		.clk        (clk_clk),                                    //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),        // reset.reset_n
		.address    (mm_interconnect_0_tt_timer_1_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_tt_timer_1_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_tt_timer_1_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_tt_timer_1_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_tt_timer_1_s1_write),     //      .write_n
		.irq        (irq_mapper_001_receiver0_irq)                //   irq.irq
	);

	slave_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                               (clk_clk),                                                     //                             clk_0_clk.clk
		.ET_Core_reset_n_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                          // ET_Core_reset_n_reset_bridge_in_reset.reset
		.ET_Core_data_master_address                 (et_core_data_master_address),                                 //                   ET_Core_data_master.address
		.ET_Core_data_master_waitrequest             (et_core_data_master_waitrequest),                             //                                      .waitrequest
		.ET_Core_data_master_byteenable              (et_core_data_master_byteenable),                              //                                      .byteenable
		.ET_Core_data_master_read                    (et_core_data_master_read),                                    //                                      .read
		.ET_Core_data_master_readdata                (et_core_data_master_readdata),                                //                                      .readdata
		.ET_Core_data_master_write                   (et_core_data_master_write),                                   //                                      .write
		.ET_Core_data_master_writedata               (et_core_data_master_writedata),                               //                                      .writedata
		.ET_Core_data_master_debugaccess             (et_core_data_master_debugaccess),                             //                                      .debugaccess
		.ET_Core_instruction_master_address          (et_core_instruction_master_address),                          //            ET_Core_instruction_master.address
		.ET_Core_instruction_master_waitrequest      (et_core_instruction_master_waitrequest),                      //                                      .waitrequest
		.ET_Core_instruction_master_read             (et_core_instruction_master_read),                             //                                      .read
		.ET_Core_instruction_master_readdata         (et_core_instruction_master_readdata),                         //                                      .readdata
		.TT_Core_data_master_address                 (tt_core_data_master_address),                                 //                   TT_Core_data_master.address
		.TT_Core_data_master_waitrequest             (tt_core_data_master_waitrequest),                             //                                      .waitrequest
		.TT_Core_data_master_byteenable              (tt_core_data_master_byteenable),                              //                                      .byteenable
		.TT_Core_data_master_read                    (tt_core_data_master_read),                                    //                                      .read
		.TT_Core_data_master_readdata                (tt_core_data_master_readdata),                                //                                      .readdata
		.TT_Core_data_master_write                   (tt_core_data_master_write),                                   //                                      .write
		.TT_Core_data_master_writedata               (tt_core_data_master_writedata),                               //                                      .writedata
		.TT_Core_data_master_debugaccess             (tt_core_data_master_debugaccess),                             //                                      .debugaccess
		.TT_Core_instruction_master_address          (tt_core_instruction_master_address),                          //            TT_Core_instruction_master.address
		.TT_Core_instruction_master_waitrequest      (tt_core_instruction_master_waitrequest),                      //                                      .waitrequest
		.TT_Core_instruction_master_read             (tt_core_instruction_master_read),                             //                                      .read
		.TT_Core_instruction_master_readdata         (tt_core_instruction_master_readdata),                         //                                      .readdata
		.ET_Core_jtag_debug_module_address           (mm_interconnect_0_et_core_jtag_debug_module_address),         //             ET_Core_jtag_debug_module.address
		.ET_Core_jtag_debug_module_write             (mm_interconnect_0_et_core_jtag_debug_module_write),           //                                      .write
		.ET_Core_jtag_debug_module_read              (mm_interconnect_0_et_core_jtag_debug_module_read),            //                                      .read
		.ET_Core_jtag_debug_module_readdata          (mm_interconnect_0_et_core_jtag_debug_module_readdata),        //                                      .readdata
		.ET_Core_jtag_debug_module_writedata         (mm_interconnect_0_et_core_jtag_debug_module_writedata),       //                                      .writedata
		.ET_Core_jtag_debug_module_byteenable        (mm_interconnect_0_et_core_jtag_debug_module_byteenable),      //                                      .byteenable
		.ET_Core_jtag_debug_module_waitrequest       (mm_interconnect_0_et_core_jtag_debug_module_waitrequest),     //                                      .waitrequest
		.ET_Core_jtag_debug_module_debugaccess       (mm_interconnect_0_et_core_jtag_debug_module_debugaccess),     //                                      .debugaccess
		.ET_Core_Memory_s1_address                   (mm_interconnect_0_et_core_memory_s1_address),                 //                     ET_Core_Memory_s1.address
		.ET_Core_Memory_s1_write                     (mm_interconnect_0_et_core_memory_s1_write),                   //                                      .write
		.ET_Core_Memory_s1_readdata                  (mm_interconnect_0_et_core_memory_s1_readdata),                //                                      .readdata
		.ET_Core_Memory_s1_writedata                 (mm_interconnect_0_et_core_memory_s1_writedata),               //                                      .writedata
		.ET_Core_Memory_s1_byteenable                (mm_interconnect_0_et_core_memory_s1_byteenable),              //                                      .byteenable
		.ET_Core_Memory_s1_chipselect                (mm_interconnect_0_et_core_memory_s1_chipselect),              //                                      .chipselect
		.ET_Core_Memory_s1_clken                     (mm_interconnect_0_et_core_memory_s1_clken),                   //                                      .clken
		.et_leds1_s1_address                         (mm_interconnect_0_et_leds1_s1_address),                       //                           et_leds1_s1.address
		.et_leds1_s1_write                           (mm_interconnect_0_et_leds1_s1_write),                         //                                      .write
		.et_leds1_s1_readdata                        (mm_interconnect_0_et_leds1_s1_readdata),                      //                                      .readdata
		.et_leds1_s1_writedata                       (mm_interconnect_0_et_leds1_s1_writedata),                     //                                      .writedata
		.et_leds1_s1_chipselect                      (mm_interconnect_0_et_leds1_s1_chipselect),                    //                                      .chipselect
		.et_leds2_s1_address                         (mm_interconnect_0_et_leds2_s1_address),                       //                           et_leds2_s1.address
		.et_leds2_s1_write                           (mm_interconnect_0_et_leds2_s1_write),                         //                                      .write
		.et_leds2_s1_readdata                        (mm_interconnect_0_et_leds2_s1_readdata),                      //                                      .readdata
		.et_leds2_s1_writedata                       (mm_interconnect_0_et_leds2_s1_writedata),                     //                                      .writedata
		.et_leds2_s1_chipselect                      (mm_interconnect_0_et_leds2_s1_chipselect),                    //                                      .chipselect
		.et_pb_1_s1_address                          (mm_interconnect_0_et_pb_1_s1_address),                        //                            et_pb_1_s1.address
		.et_pb_1_s1_readdata                         (mm_interconnect_0_et_pb_1_s1_readdata),                       //                                      .readdata
		.et_pb_2_s1_address                          (mm_interconnect_0_et_pb_2_s1_address),                        //                            et_pb_2_s1.address
		.et_pb_2_s1_readdata                         (mm_interconnect_0_et_pb_2_s1_readdata),                       //                                      .readdata
		.et_spi_0_spi_control_port_address           (mm_interconnect_0_et_spi_0_spi_control_port_address),         //             et_spi_0_spi_control_port.address
		.et_spi_0_spi_control_port_write             (mm_interconnect_0_et_spi_0_spi_control_port_write),           //                                      .write
		.et_spi_0_spi_control_port_read              (mm_interconnect_0_et_spi_0_spi_control_port_read),            //                                      .read
		.et_spi_0_spi_control_port_readdata          (mm_interconnect_0_et_spi_0_spi_control_port_readdata),        //                                      .readdata
		.et_spi_0_spi_control_port_writedata         (mm_interconnect_0_et_spi_0_spi_control_port_writedata),       //                                      .writedata
		.et_spi_0_spi_control_port_chipselect        (mm_interconnect_0_et_spi_0_spi_control_port_chipselect),      //                                      .chipselect
		.et_spican_int_s1_address                    (mm_interconnect_0_et_spican_int_s1_address),                  //                      et_spican_int_s1.address
		.et_spican_int_s1_write                      (mm_interconnect_0_et_spican_int_s1_write),                    //                                      .write
		.et_spican_int_s1_readdata                   (mm_interconnect_0_et_spican_int_s1_readdata),                 //                                      .readdata
		.et_spican_int_s1_writedata                  (mm_interconnect_0_et_spican_int_s1_writedata),                //                                      .writedata
		.et_spican_int_s1_chipselect                 (mm_interconnect_0_et_spican_int_s1_chipselect),               //                                      .chipselect
		.jtag_uart_0_avalon_jtag_slave_address       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //         jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                      .write
		.jtag_uart_0_avalon_jtag_slave_read          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                      .read
		.jtag_uart_0_avalon_jtag_slave_readdata      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                      .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                      .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                      .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                      .chipselect
		.msg_buf_mutex_s1_address                    (mm_interconnect_0_msg_buf_mutex_s1_address),                  //                      msg_buf_mutex_s1.address
		.msg_buf_mutex_s1_write                      (mm_interconnect_0_msg_buf_mutex_s1_write),                    //                                      .write
		.msg_buf_mutex_s1_read                       (mm_interconnect_0_msg_buf_mutex_s1_read),                     //                                      .read
		.msg_buf_mutex_s1_readdata                   (mm_interconnect_0_msg_buf_mutex_s1_readdata),                 //                                      .readdata
		.msg_buf_mutex_s1_writedata                  (mm_interconnect_0_msg_buf_mutex_s1_writedata),                //                                      .writedata
		.msg_buf_mutex_s1_chipselect                 (mm_interconnect_0_msg_buf_mutex_s1_chipselect),               //                                      .chipselect
		.msg_buf_ram_s1_address                      (mm_interconnect_0_msg_buf_ram_s1_address),                    //                        msg_buf_ram_s1.address
		.msg_buf_ram_s1_write                        (mm_interconnect_0_msg_buf_ram_s1_write),                      //                                      .write
		.msg_buf_ram_s1_readdata                     (mm_interconnect_0_msg_buf_ram_s1_readdata),                   //                                      .readdata
		.msg_buf_ram_s1_writedata                    (mm_interconnect_0_msg_buf_ram_s1_writedata),                  //                                      .writedata
		.msg_buf_ram_s1_byteenable                   (mm_interconnect_0_msg_buf_ram_s1_byteenable),                 //                                      .byteenable
		.msg_buf_ram_s1_chipselect                   (mm_interconnect_0_msg_buf_ram_s1_chipselect),                 //                                      .chipselect
		.msg_buf_ram_s1_clken                        (mm_interconnect_0_msg_buf_ram_s1_clken),                      //                                      .clken
		.pio_0_s1_address                            (mm_interconnect_0_pio_0_s1_address),                          //                              pio_0_s1.address
		.pio_0_s1_write                              (mm_interconnect_0_pio_0_s1_write),                            //                                      .write
		.pio_0_s1_readdata                           (mm_interconnect_0_pio_0_s1_readdata),                         //                                      .readdata
		.pio_0_s1_writedata                          (mm_interconnect_0_pio_0_s1_writedata),                        //                                      .writedata
		.pio_0_s1_chipselect                         (mm_interconnect_0_pio_0_s1_chipselect),                       //                                      .chipselect
		.TT_Core_jtag_debug_module_address           (mm_interconnect_0_tt_core_jtag_debug_module_address),         //             TT_Core_jtag_debug_module.address
		.TT_Core_jtag_debug_module_write             (mm_interconnect_0_tt_core_jtag_debug_module_write),           //                                      .write
		.TT_Core_jtag_debug_module_read              (mm_interconnect_0_tt_core_jtag_debug_module_read),            //                                      .read
		.TT_Core_jtag_debug_module_readdata          (mm_interconnect_0_tt_core_jtag_debug_module_readdata),        //                                      .readdata
		.TT_Core_jtag_debug_module_writedata         (mm_interconnect_0_tt_core_jtag_debug_module_writedata),       //                                      .writedata
		.TT_Core_jtag_debug_module_byteenable        (mm_interconnect_0_tt_core_jtag_debug_module_byteenable),      //                                      .byteenable
		.TT_Core_jtag_debug_module_waitrequest       (mm_interconnect_0_tt_core_jtag_debug_module_waitrequest),     //                                      .waitrequest
		.TT_Core_jtag_debug_module_debugaccess       (mm_interconnect_0_tt_core_jtag_debug_module_debugaccess),     //                                      .debugaccess
		.TT_core_memory_s1_address                   (mm_interconnect_0_tt_core_memory_s1_address),                 //                     TT_core_memory_s1.address
		.TT_core_memory_s1_write                     (mm_interconnect_0_tt_core_memory_s1_write),                   //                                      .write
		.TT_core_memory_s1_readdata                  (mm_interconnect_0_tt_core_memory_s1_readdata),                //                                      .readdata
		.TT_core_memory_s1_writedata                 (mm_interconnect_0_tt_core_memory_s1_writedata),               //                                      .writedata
		.TT_core_memory_s1_byteenable                (mm_interconnect_0_tt_core_memory_s1_byteenable),              //                                      .byteenable
		.TT_core_memory_s1_chipselect                (mm_interconnect_0_tt_core_memory_s1_chipselect),              //                                      .chipselect
		.TT_core_memory_s1_clken                     (mm_interconnect_0_tt_core_memory_s1_clken),                   //                                      .clken
		.tt_leds_s1_address                          (mm_interconnect_0_tt_leds_s1_address),                        //                            tt_leds_s1.address
		.tt_leds_s1_write                            (mm_interconnect_0_tt_leds_s1_write),                          //                                      .write
		.tt_leds_s1_readdata                         (mm_interconnect_0_tt_leds_s1_readdata),                       //                                      .readdata
		.tt_leds_s1_writedata                        (mm_interconnect_0_tt_leds_s1_writedata),                      //                                      .writedata
		.tt_leds_s1_chipselect                       (mm_interconnect_0_tt_leds_s1_chipselect),                     //                                      .chipselect
		.tt_pb_1_s1_address                          (mm_interconnect_0_tt_pb_1_s1_address),                        //                            tt_pb_1_s1.address
		.tt_pb_1_s1_readdata                         (mm_interconnect_0_tt_pb_1_s1_readdata),                       //                                      .readdata
		.tt_timer_1_s1_address                       (mm_interconnect_0_tt_timer_1_s1_address),                     //                         tt_timer_1_s1.address
		.tt_timer_1_s1_write                         (mm_interconnect_0_tt_timer_1_s1_write),                       //                                      .write
		.tt_timer_1_s1_readdata                      (mm_interconnect_0_tt_timer_1_s1_readdata),                    //                                      .readdata
		.tt_timer_1_s1_writedata                     (mm_interconnect_0_tt_timer_1_s1_writedata),                   //                                      .writedata
		.tt_timer_1_s1_chipselect                    (mm_interconnect_0_tt_timer_1_s1_chipselect)                   //                                      .chipselect
	);

	slave_irq_mapper irq_mapper (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.sender_irq    (et_core_d_irq_irq)                   //    sender.irq
	);

	slave_irq_mapper_001 irq_mapper_001 (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_001_receiver0_irq),       // receiver0.irq
		.sender_irq    (tt_core_d_irq_irq)                   //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (tt_core_jtag_debug_module_reset_reset), // reset_in0.reset
		.reset_in1      (et_core_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (),                                      //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),        // reset_out.reset
		.reset_req      (),                                      // (terminated)
		.reset_req_in0  (1'b0),                                  // (terminated)
		.reset_req_in1  (1'b0),                                  // (terminated)
		.reset_in2      (1'b0),                                  // (terminated)
		.reset_req_in2  (1'b0),                                  // (terminated)
		.reset_in3      (1'b0),                                  // (terminated)
		.reset_req_in3  (1'b0),                                  // (terminated)
		.reset_in4      (1'b0),                                  // (terminated)
		.reset_req_in4  (1'b0),                                  // (terminated)
		.reset_in5      (1'b0),                                  // (terminated)
		.reset_req_in5  (1'b0),                                  // (terminated)
		.reset_in6      (1'b0),                                  // (terminated)
		.reset_req_in6  (1'b0),                                  // (terminated)
		.reset_in7      (1'b0),                                  // (terminated)
		.reset_req_in7  (1'b0),                                  // (terminated)
		.reset_in8      (1'b0),                                  // (terminated)
		.reset_req_in8  (1'b0),                                  // (terminated)
		.reset_in9      (1'b0),                                  // (terminated)
		.reset_req_in9  (1'b0),                                  // (terminated)
		.reset_in10     (1'b0),                                  // (terminated)
		.reset_req_in10 (1'b0),                                  // (terminated)
		.reset_in11     (1'b0),                                  // (terminated)
		.reset_req_in11 (1'b0),                                  // (terminated)
		.reset_in12     (1'b0),                                  // (terminated)
		.reset_req_in12 (1'b0),                                  // (terminated)
		.reset_in13     (1'b0),                                  // (terminated)
		.reset_req_in13 (1'b0),                                  // (terminated)
		.reset_in14     (1'b0),                                  // (terminated)
		.reset_req_in14 (1'b0),                                  // (terminated)
		.reset_in15     (1'b0),                                  // (terminated)
		.reset_req_in15 (1'b0)                                   // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (rst_controller_reset_out_reset),         // reset_in0.reset
		.reset_in1      (et_core_jtag_debug_module_reset_reset),  // reset_in1.reset
		.reset_in2      (tt_core_jtag_debug_module_reset_reset),  // reset_in2.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
